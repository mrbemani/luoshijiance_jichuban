/**
 * Web server for web access and api call.
 */


module webserver

import math



